library verilog;
use verilog.vl_types.all;
entity lab5_test is
end lab5_test;
