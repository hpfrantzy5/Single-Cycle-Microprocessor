`ifndef _LAB_5_IRAM_V_
`define _LAB_5_IRAM_V_

module lab5iram
(
  input         CLK,
  input         RESET,
  input  [ 7:0] ADDR,
  output [15:0] Q
);

  reg  [15:0] mem [0:127]; // Instruction memory with 16 bit entries.
  wire [ 6:0] SADDR;
  integer     i;

  assign SADDR = ADDR[7:1];
  assign Q     = mem[SADDR];

  always @ ( posedge CLK )
  begin
    if ( RESET ) begin
         mem[0]  <= 16'b1111010010010001; //SUB  R2, R2,    R2
         mem[1]  <= 16'b1111001001001001; //SUB  R1, R1,    R1
         mem[2]  <= 16'b0101010010111111; //ADDI R2, R2,    -1
         mem[3]  <= 16'b0101010010111111; //ADDI R2, R2,    -1
         mem[4]  <= 16'b0101010010111111; //ADDI R2, R2,    -1
         mem[5]  <= 16'b0101010010111111; //ADDI R2, R2,    -1
         mem[6]  <= 16'b0101010010000011; //ADDI R2, R2,     3
         mem[7]  <= 16'b0100010001000000; //SB   R1, 0(R2)
         mem[8]  <= 16'b0101001001000001; //ADDI R1, R1,     1
         mem[9]  <= 16'b0100010001000000; //SB   R1, 0(R2)
         mem[10] <= 16'b0101001001000001; //ADDI R1, R1,     1
         mem[11] <= 16'b0100010001000000; //SB   R1, 0(R2)
         mem[12] <= 16'b0101001001000001; //ADDI R1, R1,     1
         mem[13] <= 16'b0100010001000000; //SB   R1, 0(R2)
         mem[14] <= 16'b0101001001000001; //ADDI R1, R1,     1
         mem[15] <= 16'b0100010001000000; //SB   R1, 0(R2)
         mem[16] <= 16'b0101001001000001; //ADDI R1, R1,     1
         mem[17] <= 16'b0100010001000000; //SB   R1, 0(R2)

         for(i = 18; i < 128; i = i + 1)
            mem[i] <= 16'b0000000000000000;
      end
  end

endmodule

`endif /* _LAB_5_IRAM_V_ */